-- Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.27.11:20:48

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module is
	port (
		data_out  : out std_logic_vector(23 downto 0);                    --  data_out.wire
		write     : in  std_logic                     := '0';             --     write.wire
		writedata : in  std_logic_vector(31 downto 0) := (others => '0'); -- writedata.wire
		data_in   : in  std_logic_vector(23 downto 0) := (others => '0'); --   data_in.wire
		sop       : in  std_logic                     := '0';             --       sop.wire
		addr      : in  std_logic_vector(1 downto 0)  := (others => '0'); --      addr.wire
		eop       : in  std_logic                     := '0';             --       eop.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0'              --          .reset
	);
end entity Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module;

architecture rtl of Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNLF52SJQ3 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNLF52SJQ3;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_multiplexer_GNCALBUTDR is
		generic (
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0;
			width                  : positive := 8;
			pipeline               : natural  := 0;
			number_inputs          : natural  := 4
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(23 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNCALBUTDR;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Binarization_Module is
		port (
			data_out : out std_logic_vector(23 downto 0);                    -- wire
			data_in  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			Clock    : in  std_logic                     := 'X';             -- clk
			aclr     : in  std_logic                     := 'X';             -- reset
			thr      : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- wire
		);
	end component Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Binarization_Module;

	component alt_dspbuilder_constant_GNZEH3JAKA is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNZEH3JAKA;

	component alt_dspbuilder_port_GN6TDLHAW6 is
		port (
			input  : in  std_logic_vector(1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN6TDLHAW6;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_constant_GNNKZSYI73 is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNNKZSYI73;

	component alt_dspbuilder_delay_GNUECIBFDH is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNUECIBFDH;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_decoder_GNM4LOIHXZ is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNM4LOIHXZ;

	component alt_dspbuilder_decoder_GNSCEXJCJK is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNSCEXJCJK;

	component alt_dspbuilder_delay_GNHYCSAEGT is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNHYCSAEGT;

	component alt_dspbuilder_delay_GNVTJPHWYT is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNVTJPHWYT;

	component alt_dspbuilder_if_statement_GN7VA7SRUP is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			c    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GN7VA7SRUP;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Gray_Module is
		port (
			Clock    : in  std_logic                     := 'X';             -- clk
			aclr     : in  std_logic                     := 'X';             -- reset
			data_in  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			data_out : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Gray_Module;

	component alt_dspbuilder_decoder_GNEQGKKPXW is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNEQGKKPXW;

	component alt_dspbuilder_cast_GNZ5LMFB5D is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(0 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNZ5LMFB5D;

	component alt_dspbuilder_cast_GNSB3OXIQS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                        -- wire
		);
	end component alt_dspbuilder_cast_GNSB3OXIQS;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	signal multiplexeruser_aclrgnd_output_wire                                            : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire                                                  : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal decoder2sclrgnd_output_wire                                                    : std_logic;                     -- Decoder2sclrGND:output -> Decoder2:sclr
	signal decoder2enavcc_output_wire                                                     : std_logic;                     -- Decoder2enaVCC:output -> Decoder2:ena
	signal decoder3sclrgnd_output_wire                                                    : std_logic;                     -- Decoder3sclrGND:output -> Decoder3:sclr
	signal decoder3enavcc_output_wire                                                     : std_logic;                     -- Decoder3enaVCC:output -> Decoder3:ena
	signal decoder1sclrgnd_output_wire                                                    : std_logic;                     -- Decoder1sclrGND:output -> Decoder1:sclr
	signal decoder1enavcc_output_wire                                                     : std_logic;                     -- Decoder1enaVCC:output -> Decoder1:ena
	signal delay6sclrgnd_output_wire                                                      : std_logic;                     -- Delay6sclrGND:output -> Delay6:sclr
	signal delay5sclrgnd_output_wire                                                      : std_logic;                     -- Delay5sclrGND:output -> Delay5:sclr
	signal delay4sclrgnd_output_wire                                                      : std_logic;                     -- Delay4sclrGND:output -> Delay4:sclr
	signal delay4enavcc_output_wire                                                       : std_logic;                     -- Delay4enaVCC:output -> Delay4:ena
	signal delay3sclrgnd_output_wire                                                      : std_logic;                     -- Delay3sclrGND:output -> Delay3:sclr
	signal delay1sclrgnd_output_wire                                                      : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal delay1enavcc_output_wire                                                       : std_logic;                     -- Delay1enaVCC:output -> Delay1:ena
	signal multiplexer2user_aclrgnd_output_wire                                           : std_logic;                     -- Multiplexer2user_aclrGND:output -> Multiplexer2:user_aclr
	signal multiplexer2enavcc_output_wire                                                 : std_logic;                     -- Multiplexer2enaVCC:output -> Multiplexer2:ena
	signal delay2sclrgnd_output_wire                                                      : std_logic;                     -- Delay2sclrGND:output -> Delay2:sclr
	signal decodersclrgnd_output_wire                                                     : std_logic;                     -- DecodersclrGND:output -> Decoder:sclr
	signal decoderenavcc_output_wire                                                      : std_logic;                     -- DecoderenaVCC:output -> Decoder:ena
	signal writedata_0_output_wire                                                        : std_logic_vector(31 downto 0); -- writedata_0:output -> [Bus_Conversion1:input, Bus_Conversion6:input]
	signal addr_0_output_wire                                                             : std_logic_vector(1 downto 0);  -- addr_0:output -> [Decoder2:data, Decoder:data]
	signal bus_conversion1_output_wire                                                    : std_logic_vector(7 downto 0);  -- Bus_Conversion1:output -> Delay2:input
	signal delay2_output_wire                                                             : std_logic_vector(7 downto 0);  -- Delay2:output -> Delay3:input
	signal delay3_output_wire                                                             : std_logic_vector(7 downto 0);  -- Delay3:output -> Gray_Binarization_Gray_Binarization_Module_Binarization_Module_0:thr
	signal delay4_output_wire                                                             : std_logic_vector(0 downto 0);  -- Delay4:output -> [Delay:input, cast2:input]
	signal bus_conversion6_output_wire                                                    : std_logic_vector(0 downto 0);  -- Bus_Conversion6:output -> Delay5:input
	signal delay5_output_wire                                                             : std_logic_vector(0 downto 0);  -- Delay5:output -> Delay6:input
	signal data_in_0_output_wire                                                          : std_logic_vector(23 downto 0); -- data_in_0:output -> [Decoder1:data, Decoder3:data, Gray_Binarization_Gray_Binarization_Module_Gray_Module_0:data_in, If_Statement1:a, Multiplexer:in0]
	signal gray_binarization_gray_binarization_module_gray_module_0_data_out_wire         : std_logic_vector(23 downto 0); -- Gray_Binarization_Gray_Binarization_Module_Gray_Module_0:data_out -> [Gray_Binarization_Gray_Binarization_Module_Binarization_Module_0:data_in, Multiplexer2:in0]
	signal constant3_output_wire                                                          : std_logic_vector(23 downto 0); -- Constant3:output -> If_Statement1:b
	signal constant4_output_wire                                                          : std_logic_vector(23 downto 0); -- Constant4:output -> If_Statement1:c
	signal if_statement1_true_wire                                                        : std_logic;                     -- If_Statement1:true -> Logical_Bit_Operator:data0
	signal sop_0_output_wire                                                              : std_logic;                     -- sop_0:output -> [Logical_Bit_Operator3:data0, Logical_Bit_Operator5:data0, Logical_Bit_Operator:data1]
	signal eop_0_output_wire                                                              : std_logic;                     -- eop_0:output -> Logical_Bit_Operator1:data0
	signal decoder_dec_wire                                                               : std_logic;                     -- Decoder:dec -> Logical_Bit_Operator2:data0
	signal write_0_output_wire                                                            : std_logic;                     -- write_0:output -> [Logical_Bit_Operator2:data1, Logical_Bit_Operator4:data1]
	signal logical_bit_operator2_result_wire                                              : std_logic;                     -- Logical_Bit_Operator2:result -> Delay2:ena
	signal decoder1_dec_wire                                                              : std_logic;                     -- Decoder1:dec -> Logical_Bit_Operator3:data1
	signal logical_bit_operator3_result_wire                                              : std_logic;                     -- Logical_Bit_Operator3:result -> Delay3:ena
	signal decoder2_dec_wire                                                              : std_logic;                     -- Decoder2:dec -> Logical_Bit_Operator4:data0
	signal logical_bit_operator4_result_wire                                              : std_logic;                     -- Logical_Bit_Operator4:result -> Delay5:ena
	signal decoder3_dec_wire                                                              : std_logic;                     -- Decoder3:dec -> Logical_Bit_Operator5:data1
	signal logical_bit_operator5_result_wire                                              : std_logic;                     -- Logical_Bit_Operator5:result -> Delay6:ena
	signal delay_output_wire                                                              : std_logic_vector(0 downto 0);  -- Delay:output -> [Multiplexer:sel, cast4:input]
	signal delay6_output_wire                                                             : std_logic_vector(0 downto 0);  -- Delay6:output -> Multiplexer2:sel
	signal gray_binarization_gray_binarization_module_binarization_module_0_data_out_wire : std_logic_vector(23 downto 0); -- Gray_Binarization_Gray_Binarization_Module_Binarization_Module_0:data_out -> Multiplexer2:in1
	signal multiplexer2_result_wire                                                       : std_logic_vector(23 downto 0); -- Multiplexer2:result -> Multiplexer:in1
	signal multiplexer_result_wire                                                        : std_logic_vector(23 downto 0); -- Multiplexer:result -> data_out_0:input
	signal delay1_output_wire                                                             : std_logic_vector(0 downto 0);  -- Delay1:output -> cast1:input
	signal cast1_output_wire                                                              : std_logic;                     -- cast1:output -> Delay:sclr
	signal cast2_output_wire                                                              : std_logic;                     -- cast2:output -> Delay:ena
	signal logical_bit_operator_result_wire                                               : std_logic;                     -- Logical_Bit_Operator:result -> cast3:input
	signal cast3_output_wire                                                              : std_logic_vector(0 downto 0);  -- cast3:output -> Delay4:input
	signal cast4_output_wire                                                              : std_logic;                     -- cast4:output -> Logical_Bit_Operator1:data1
	signal logical_bit_operator1_result_wire                                              : std_logic;                     -- Logical_Bit_Operator1:result -> cast5:input
	signal cast5_output_wire                                                              : std_logic_vector(0 downto 0);  -- cast5:output -> Delay1:input
	signal clock_0_clock_output_reset                                                     : std_logic;                     -- Clock_0:aclr_out -> [Decoder1:aclr, Decoder2:aclr, Decoder3:aclr, Decoder:aclr, Delay1:aclr, Delay2:aclr, Delay3:aclr, Delay4:aclr, Delay5:aclr, Delay6:aclr, Delay:aclr, Gray_Binarization_Gray_Binarization_Module_Binarization_Module_0:aclr, Gray_Binarization_Gray_Binarization_Module_Gray_Module_0:aclr, Multiplexer2:aclr, Multiplexer:aclr]
	signal clock_0_clock_output_clk                                                       : std_logic;                     -- Clock_0:clock_out -> [Decoder1:clock, Decoder2:clock, Decoder3:clock, Decoder:clock, Delay1:clock, Delay2:clock, Delay3:clock, Delay4:clock, Delay5:clock, Delay6:clock, Delay:clock, Gray_Binarization_Gray_Binarization_Module_Binarization_Module_0:Clock, Gray_Binarization_Gray_Binarization_Module_Gray_Module_0:Clock, Multiplexer2:clock, Multiplexer:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion1 : component alt_dspbuilder_cast_GNLF52SJQ3
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => writedata_0_output_wire,     --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	writedata_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => writedata,               --  input.wire
			output => writedata_0_output_wire  -- output.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNCALBUTDR
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0,
			width                  => 24,
			pipeline               => 0,
			number_inputs          => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => delay_output_wire,                   --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => data_in_0_output_wire,               --        in0.wire
			in1       => multiplexer2_result_wire             --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	gray_binarization_gray_binarization_module_binarization_module_0 : component Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Binarization_Module
		port map (
			data_out => gray_binarization_gray_binarization_module_binarization_module_0_data_out_wire, -- data_out.wire
			data_in  => gray_binarization_gray_binarization_module_gray_module_0_data_out_wire,         --  data_in.wire
			Clock    => clock_0_clock_output_clk,                                                       --    Clock.clk
			aclr     => clock_0_clock_output_reset,                                                     --         .reset
			thr      => delay3_output_wire                                                              --      thr.wire
		);

	constant4 : component alt_dspbuilder_constant_GNZEH3JAKA
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000001111",
			width      => 24
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	addr_0 : component alt_dspbuilder_port_GN6TDLHAW6
		port map (
			input  => addr,               --  input.wire
			output => addr_0_output_wire  -- output.wire
		);

	logical_bit_operator5 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator5_result_wire, -- result.wire
			data0  => sop_0_output_wire,                 --  data0.wire
			data1  => decoder3_dec_wire                  --  data1.wire
		);

	logical_bit_operator4 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator4_result_wire, -- result.wire
			data0  => decoder2_dec_wire,                 --  data0.wire
			data1  => write_0_output_wire                --  data1.wire
		);

	constant3 : component alt_dspbuilder_constant_GNNKZSYI73
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	delay : component alt_dspbuilder_delay_GNUECIBFDH
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => delay4_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay_output_wire,          --     output.wire
			sclr   => cast1_output_wire,          --       sclr.wire
			ena    => cast2_output_wire           --        ena.wire
		);

	write_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => write,               --  input.wire
			output => write_0_output_wire  -- output.wire
		);

	logical_bit_operator3 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator3_result_wire, -- result.wire
			data0  => sop_0_output_wire,                 --  data0.wire
			data1  => decoder1_dec_wire                  --  data1.wire
		);

	logical_bit_operator2 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator2_result_wire, -- result.wire
			data0  => decoder_dec_wire,                  --  data0.wire
			data1  => write_0_output_wire                --  data1.wire
		);

	eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eop,               --  input.wire
			output => eop_0_output_wire  -- output.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire, -- result.wire
			data0  => eop_0_output_wire,                 --  data0.wire
			data1  => cast4_output_wire                  --  data1.wire
		);

	decoder2 : component alt_dspbuilder_decoder_GNM4LOIHXZ
		generic map (
			decode   => "01",
			pipeline => 1,
			width    => 2
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => addr_0_output_wire,          --       data.wire
			dec   => decoder2_dec_wire,           --        dec.wire
			sclr  => decoder2sclrgnd_output_wire, --       sclr.wire
			ena   => decoder2enavcc_output_wire   --        ena.wire
		);

	decoder2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder2sclrgnd_output_wire  -- output.wire
		);

	decoder2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder2enavcc_output_wire  -- output.wire
		);

	decoder3 : component alt_dspbuilder_decoder_GNSCEXJCJK
		generic map (
			decode   => "000000000000000000001111",
			pipeline => 0,
			width    => 24
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => data_in_0_output_wire,       --       data.wire
			dec   => decoder3_dec_wire,           --        dec.wire
			sclr  => decoder3sclrgnd_output_wire, --       sclr.wire
			ena   => decoder3enavcc_output_wire   --        ena.wire
		);

	decoder3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder3sclrgnd_output_wire  -- output.wire
		);

	decoder3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder3enavcc_output_wire  -- output.wire
		);

	decoder1 : component alt_dspbuilder_decoder_GNSCEXJCJK
		generic map (
			decode   => "000000000000000000001111",
			pipeline => 0,
			width    => 24
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => data_in_0_output_wire,       --       data.wire
			dec   => decoder1_dec_wire,           --        dec.wire
			sclr  => decoder1sclrgnd_output_wire, --       sclr.wire
			ena   => decoder1enavcc_output_wire   --        ena.wire
		);

	decoder1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder1sclrgnd_output_wire  -- output.wire
		);

	decoder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder1enavcc_output_wire  -- output.wire
		);

	logical_bit_operator : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator_result_wire, -- result.wire
			data0  => if_statement1_true_wire,          --  data0.wire
			data1  => sop_0_output_wire                 --  data1.wire
		);

	delay6 : component alt_dspbuilder_delay_GNUECIBFDH
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => delay5_output_wire,                --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay6_output_wire,                --     output.wire
			sclr   => delay6sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator5_result_wire  --        ena.wire
		);

	delay6sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay6sclrgnd_output_wire  -- output.wire
		);

	delay5 : component alt_dspbuilder_delay_GNUECIBFDH
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => bus_conversion6_output_wire,       --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay5_output_wire,                --     output.wire
			sclr   => delay5sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator4_result_wire  --        ena.wire
		);

	delay5sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay5sclrgnd_output_wire  -- output.wire
		);

	delay4 : component alt_dspbuilder_delay_GNHYCSAEGT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => cast3_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay4_output_wire,         --     output.wire
			sclr   => delay4sclrgnd_output_wire,  --       sclr.wire
			ena    => delay4enavcc_output_wire    --        ena.wire
		);

	delay4sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay4sclrgnd_output_wire  -- output.wire
		);

	delay4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay4enavcc_output_wire  -- output.wire
		);

	delay3 : component alt_dspbuilder_delay_GNVTJPHWYT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "01111111",
			width      => 8
		)
		port map (
			input  => delay2_output_wire,                --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay3_output_wire,                --     output.wire
			sclr   => delay3sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator3_result_wire  --        ena.wire
		);

	delay3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay3sclrgnd_output_wire  -- output.wire
		);

	if_statement1 : component alt_dspbuilder_if_statement_GN7VA7SRUP
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(a=b) and (a /= c)",
			number_inputs   => 3,
			width           => 24
		)
		port map (
			true => if_statement1_true_wire, -- true.wire
			a    => data_in_0_output_wire,   --    a.wire
			b    => constant3_output_wire,   --    b.wire
			c    => constant4_output_wire    --    c.wire
		);

	sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sop,               --  input.wire
			output => sop_0_output_wire  -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNHYCSAEGT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => cast5_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay1_output_wire,         --     output.wire
			sclr   => delay1sclrgnd_output_wire,  --       sclr.wire
			ena    => delay1enavcc_output_wire    --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	delay1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay1enavcc_output_wire  -- output.wire
		);

	multiplexer2 : component alt_dspbuilder_multiplexer_GNCALBUTDR
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0,
			width                  => 24,
			pipeline               => 0,
			number_inputs          => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,                                                       -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                                     --           .reset
			sel       => delay6_output_wire,                                                             --        sel.wire
			result    => multiplexer2_result_wire,                                                       --     result.wire
			ena       => multiplexer2enavcc_output_wire,                                                 --        ena.wire
			user_aclr => multiplexer2user_aclrgnd_output_wire,                                           --  user_aclr.wire
			in0       => gray_binarization_gray_binarization_module_gray_module_0_data_out_wire,         --        in0.wire
			in1       => gray_binarization_gray_binarization_module_binarization_module_0_data_out_wire  --        in1.wire
		);

	multiplexer2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer2user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer2enavcc_output_wire  -- output.wire
		);

	delay2 : component alt_dspbuilder_delay_GNVTJPHWYT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "01111111",
			width      => 8
		)
		port map (
			input  => bus_conversion1_output_wire,       --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay2_output_wire,                --     output.wire
			sclr   => delay2sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator2_result_wire  --        ena.wire
		);

	delay2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay2sclrgnd_output_wire  -- output.wire
		);

	data_out_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => data_out                 -- output.wire
		);

	gray_binarization_gray_binarization_module_gray_module_0 : component Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Gray_Module
		port map (
			Clock    => clock_0_clock_output_clk,                                               --    Clock.clk
			aclr     => clock_0_clock_output_reset,                                             --         .reset
			data_in  => data_in_0_output_wire,                                                  --  data_in.wire
			data_out => gray_binarization_gray_binarization_module_gray_module_0_data_out_wire  -- data_out.wire
		);

	data_in_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => data_in,               --  input.wire
			output => data_in_0_output_wire  -- output.wire
		);

	decoder : component alt_dspbuilder_decoder_GNEQGKKPXW
		generic map (
			decode   => "10",
			pipeline => 1,
			width    => 2
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			data  => addr_0_output_wire,         --       data.wire
			dec   => decoder_dec_wire,           --        dec.wire
			sclr  => decodersclrgnd_output_wire, --       sclr.wire
			ena   => decoderenavcc_output_wire   --        ena.wire
		);

	decodersclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decodersclrgnd_output_wire  -- output.wire
		);

	decoderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoderenavcc_output_wire  -- output.wire
		);

	bus_conversion6 : component alt_dspbuilder_cast_GNZ5LMFB5D
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => writedata_0_output_wire,     --  input.wire
			output => bus_conversion6_output_wire  -- output.wire
		);

	cast1 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire, --  input.wire
			output => cast1_output_wire   -- output.wire
		);

	cast2 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay4_output_wire, --  input.wire
			output => cast2_output_wire   -- output.wire
		);

	cast3 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator_result_wire, --  input.wire
			output => cast3_output_wire                 -- output.wire
		);

	cast4 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay_output_wire, --  input.wire
			output => cast4_output_wire  -- output.wire
		);

	cast5 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator1_result_wire, --  input.wire
			output => cast5_output_wire                  -- output.wire
		);

end architecture rtl; -- of Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module
