-- Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Gray_Module.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.27.11:20:48

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Gray_Module is
	port (
		Clock    : in  std_logic                     := '0';             --    Clock.clk
		aclr     : in  std_logic                     := '0';             --         .reset
		data_in  : in  std_logic_vector(23 downto 0) := (others => '0'); --  data_in.wire
		data_out : out std_logic_vector(23 downto 0)                     -- data_out.wire
	);
end entity Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Gray_Module;

architecture rtl of Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Gray_Module is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNJGR7GQ2L is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNJGR7GQ2L;

	component alt_dspbuilder_cast_GNKXX25S2S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNKXX25S2S;

	component alt_dspbuilder_cast_GN6OMCQQS7 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GN6OMCQQS7;

	component alt_dspbuilder_bus_concat_GNIIOZRPJD is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNIIOZRPJD;

	component alt_dspbuilder_barrelshifter_GNV5DVAGHT is
		generic (
			DISTANCE_WIDTH          : natural := 3;
			NDIRECTION              : natural := 0;
			SIGNED                  : integer := 1;
			use_dedicated_circuitry : string  := "false";
			PIPELINE                : natural := 0;
			WIDTH                   : natural := 8
		);
		port (
			a         : in  std_logic_vector(WIDTH-1 downto 0)          := (others => 'X'); -- wire
			aclr      : in  std_logic                                   := 'X';             -- clk
			clock     : in  std_logic                                   := 'X';             -- clk
			direction : in  std_logic                                   := 'X';             -- wire
			distance  : in  std_logic_vector(DISTANCE_WIDTH-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                                   := 'X';             -- wire
			r         : out std_logic_vector(WIDTH-1 downto 0);                             -- wire
			user_aclr : in  std_logic                                   := 'X'              -- wire
		);
	end component alt_dspbuilder_barrelshifter_GNV5DVAGHT;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_multiply_add_GNKLXFKAO3 is
		generic (
			family                  : string  := "Stratix";
			direction               : string  := "AddAdd";
			data3b_const            : string  := "00000000";
			data2b_const            : string  := "00000000";
			representation          : string  := "SIGNED";
			dataWidth               : integer := 8;
			data4b_const            : string  := "00000000";
			number_multipliers      : integer := 2;
			pipeline_register       : string  := "NoRegister";
			use_dedicated_circuitry : integer := 0;
			data1b_const            : string  := "00000000";
			use_b_consts            : natural := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			data1a    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			data2a    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			data3a    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(17 downto 0);                    -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			ena       : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_multiply_add_GNKLXFKAO3;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_constant_GNPXZ5JSVR is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(3 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNPXZ5JSVR;

	component alt_dspbuilder_bus_concat_GN55ETJ4VI is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GN55ETJ4VI;

	component alt_dspbuilder_cast_GN7IAAYCSZ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GN7IAAYCSZ;

	signal barrel_shifteruser_aclrgnd_output_wire : std_logic;                     -- Barrel_Shifteruser_aclrGND:output -> Barrel_Shifter:user_aclr
	signal barrel_shifterenavcc_output_wire       : std_logic;                     -- Barrel_ShifterenaVCC:output -> Barrel_Shifter:ena
	signal multiply_adduser_aclrgnd_output_wire   : std_logic;                     -- Multiply_Adduser_aclrGND:output -> Multiply_Add:user_aclr
	signal multiply_addenavcc_output_wire         : std_logic;                     -- Multiply_AddenaVCC:output -> Multiply_Add:ena
	signal bus_concatenation_output_wire          : std_logic_vector(15 downto 0); -- Bus_Concatenation:output -> Bus_Concatenation1:b
	signal barrel_shifter_r_wire                  : std_logic_vector(17 downto 0); -- Barrel_Shifter:r -> Bus_Conversion2:input
	signal bus_conversion2_output_wire            : std_logic_vector(7 downto 0);  -- Bus_Conversion2:output -> [Bus_Concatenation1:a, Bus_Concatenation:a, Bus_Concatenation:b]
	signal data_in_0_output_wire                  : std_logic_vector(23 downto 0); -- data_in_0:output -> [Bus_Conversion3:input, Bus_Conversion4:input, Bus_Conversion5:input]
	signal constant5_output_wire                  : std_logic_vector(3 downto 0);  -- Constant5:output -> Barrel_Shifter:distance
	signal bus_conversion5_output_wire            : std_logic_vector(7 downto 0);  -- Bus_Conversion5:output -> Multiply_Add:data1a
	signal bus_conversion4_output_wire            : std_logic_vector(7 downto 0);  -- Bus_Conversion4:output -> Multiply_Add:data2a
	signal bus_conversion3_output_wire            : std_logic_vector(7 downto 0);  -- Bus_Conversion3:output -> Multiply_Add:data3a
	signal multiply_add_result_wire               : std_logic_vector(17 downto 0); -- Multiply_Add:result -> Barrel_Shifter:a
	signal bus_concatenation1_output_wire         : std_logic_vector(23 downto 0); -- Bus_Concatenation1:output -> data_out_0:input
	signal clock_0_clock_output_reset             : std_logic;                     -- Clock_0:aclr_out -> [Barrel_Shifter:aclr, Bus_Concatenation1:aclr, Bus_Concatenation:aclr, Multiply_Add:aclr]
	signal clock_0_clock_output_clk               : std_logic;                     -- Clock_0:clock_out -> [Barrel_Shifter:clock, Bus_Concatenation1:clock, Bus_Concatenation:clock, Multiply_Add:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion2 : component alt_dspbuilder_cast_GNJGR7GQ2L
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => barrel_shifter_r_wire,       --  input.wire
			output => bus_conversion2_output_wire  -- output.wire
		);

	bus_conversion3 : component alt_dspbuilder_cast_GNKXX25S2S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_in_0_output_wire,       --  input.wire
			output => bus_conversion3_output_wire  -- output.wire
		);

	bus_conversion4 : component alt_dspbuilder_cast_GN6OMCQQS7
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_in_0_output_wire,       --  input.wire
			output => bus_conversion4_output_wire  -- output.wire
		);

	bus_concatenation : component alt_dspbuilder_bus_concat_GNIIOZRPJD
		generic map (
			widthB => 8,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,    --           .reset
			a      => bus_conversion2_output_wire,   --          a.wire
			b      => bus_conversion2_output_wire,   --          b.wire
			output => bus_concatenation_output_wire  --     output.wire
		);

	barrel_shifter : component alt_dspbuilder_barrelshifter_GNV5DVAGHT
		generic map (
			DISTANCE_WIDTH          => 4,
			NDIRECTION              => 1,
			SIGNED                  => 0,
			use_dedicated_circuitry => "false",
			PIPELINE                => 0,
			WIDTH                   => 18
		)
		port map (
			clock     => clock_0_clock_output_clk,               -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,             --           .reset
			a         => multiply_add_result_wire,               --          a.wire
			r         => barrel_shifter_r_wire,                  --          r.wire
			distance  => constant5_output_wire,                  --   distance.wire
			ena       => barrel_shifterenavcc_output_wire,       --        ena.wire
			user_aclr => barrel_shifteruser_aclrgnd_output_wire  --  user_aclr.wire
		);

	barrel_shifteruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => barrel_shifteruser_aclrgnd_output_wire  -- output.wire
		);

	barrel_shifterenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => barrel_shifterenavcc_output_wire  -- output.wire
		);

	multiply_add : component alt_dspbuilder_multiply_add_GNKLXFKAO3
		generic map (
			family                  => "Cyclone V",
			direction               => "AddAdd",
			data3b_const            => "00011110",
			data2b_const            => "10010110",
			representation          => "UNSIGNED",
			dataWidth               => 8,
			data4b_const            => "01001100",
			number_multipliers      => 3,
			pipeline_register       => "NoRegister",
			use_dedicated_circuitry => 1,
			data1b_const            => "01001100",
			use_b_consts            => 1
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			data1a    => bus_conversion5_output_wire,          --     data1a.wire
			data2a    => bus_conversion4_output_wire,          --     data2a.wire
			data3a    => bus_conversion3_output_wire,          --     data3a.wire
			result    => multiply_add_result_wire,             --     result.wire
			user_aclr => multiply_adduser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => multiply_addenavcc_output_wire        --        ena.wire
		);

	multiply_adduser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiply_adduser_aclrgnd_output_wire  -- output.wire
		);

	multiply_addenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiply_addenavcc_output_wire  -- output.wire
		);

	data_out_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => bus_concatenation1_output_wire, --  input.wire
			output => data_out                        -- output.wire
		);

	constant5 : component alt_dspbuilder_constant_GNPXZ5JSVR
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "1000",
			width      => 4
		)
		port map (
			output => constant5_output_wire  -- output.wire
		);

	data_in_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => data_in,               --  input.wire
			output => data_in_0_output_wire  -- output.wire
		);

	bus_concatenation1 : component alt_dspbuilder_bus_concat_GN55ETJ4VI
		generic map (
			widthB => 16,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_conversion2_output_wire,    --          a.wire
			b      => bus_concatenation_output_wire,  --          b.wire
			output => bus_concatenation1_output_wire  --     output.wire
		);

	bus_conversion5 : component alt_dspbuilder_cast_GN7IAAYCSZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_in_0_output_wire,       --  input.wire
			output => bus_conversion5_output_wire  -- output.wire
		);

end architecture rtl; -- of Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Gray_Module
