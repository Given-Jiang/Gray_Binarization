-- Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Binarization_Module.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.27.11:20:48

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Binarization_Module is
	port (
		data_out : out std_logic_vector(23 downto 0);                    -- data_out.wire
		data_in  : in  std_logic_vector(23 downto 0) := (others => '0'); --  data_in.wire
		Clock    : in  std_logic                     := '0';             --    Clock.clk
		aclr     : in  std_logic                     := '0';             --         .reset
		thr      : in  std_logic_vector(7 downto 0)  := (others => '0')  --      thr.wire
	);
end entity Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Binarization_Module;

architecture rtl of Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Binarization_Module is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_multiplexer_GNCALBUTDR is
		generic (
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0;
			width                  : positive := 8;
			pipeline               : natural  := 0;
			number_inputs          : natural  := 4
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(23 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNCALBUTDR;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component alt_dspbuilder_if_statement_GNYT6HZJI5 is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                       -- wire
			a    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(7 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNYT6HZJI5;

	component alt_dspbuilder_constant_GNLMV7GZFA is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNLMV7GZFA;

	component alt_dspbuilder_constant_GNNKZSYI73 is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNNKZSYI73;

	component alt_dspbuilder_cast_GNKXX25S2S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNKXX25S2S;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	signal multiplexer1user_aclrgnd_output_wire : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire       : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal data_in_0_output_wire                : std_logic_vector(23 downto 0); -- data_in_0:output -> Bus_Conversion:input
	signal bus_conversion_output_wire           : std_logic_vector(7 downto 0);  -- Bus_Conversion:output -> If_Statement:a
	signal thr_0_output_wire                    : std_logic_vector(7 downto 0);  -- thr_0:output -> If_Statement:b
	signal constant1_output_wire                : std_logic_vector(23 downto 0); -- Constant1:output -> Multiplexer1:in0
	signal constant2_output_wire                : std_logic_vector(23 downto 0); -- Constant2:output -> Multiplexer1:in1
	signal multiplexer1_result_wire             : std_logic_vector(23 downto 0); -- Multiplexer1:result -> data_out_0:input
	signal if_statement_true_wire               : std_logic;                     -- If_Statement:true -> cast0:input
	signal cast0_output_wire                    : std_logic_vector(0 downto 0);  -- cast0:output -> Multiplexer1:sel
	signal clock_0_clock_output_reset           : std_logic;                     -- Clock_0:aclr_out -> Multiplexer1:aclr
	signal clock_0_clock_output_clk             : std_logic;                     -- Clock_0:clock_out -> Multiplexer1:clock

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNCALBUTDR
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0,
			width                  => 24,
			pipeline               => 0,
			number_inputs          => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast0_output_wire,                    --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => constant1_output_wire,                --        in0.wire
			in1       => constant2_output_wire                 --        in1.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	thr_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => thr,               --  input.wire
			output => thr_0_output_wire  -- output.wire
		);

	if_statement : component alt_dspbuilder_if_statement_GNYT6HZJI5
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "a>b",
			number_inputs   => 2,
			width           => 8
		)
		port map (
			true => if_statement_true_wire,     -- true.wire
			a    => bus_conversion_output_wire, --    a.wire
			b    => thr_0_output_wire           --    b.wire
		);

	constant2 : component alt_dspbuilder_constant_GNLMV7GZFA
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "111111111111111111111111",
			width      => 24
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	constant1 : component alt_dspbuilder_constant_GNNKZSYI73
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	bus_conversion : component alt_dspbuilder_cast_GNKXX25S2S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_in_0_output_wire,      --  input.wire
			output => bus_conversion_output_wire  -- output.wire
		);

	data_out_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => multiplexer1_result_wire, --  input.wire
			output => data_out                  -- output.wire
		);

	data_in_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => data_in,               --  input.wire
			output => data_in_0_output_wire  -- output.wire
		);

	cast0 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => if_statement_true_wire, --  input.wire
			output => cast0_output_wire       -- output.wire
		);

end architecture rtl; -- of Gray_Binarization_GN_Gray_Binarization_Gray_Binarization_Module_Binarization_Module
